module assign_keyword(input [2:0] a,b,output [2:0] c);

assign c=a&b;

endmodule
